
XX1 d0 d1 d2 d3 d4 d5 d6 d7 d8 d9 N001 out 0 10bit
V1 N001 0 3.3
V2 d6 0 PULSE(0 1.8 640m 0.1p 0.1p 640m 1280m 40)
V3 d7 0 PULSE(0 1.8 1280m 0.1p 0.1p 1280m 2560m 20)
V4 d8 0 PULSE(0 1.8 2560m 0.1p 0.1p 2560m 5120m 10)
V5 d9 0 PULSE(0 1.8 5120m 0.1p 0.1p 5120m 10240m 5)
V6 d0 0 PULSE(0 1.8 10m 0.1p 0.1p 10m 20m 200)
V7 d1 0 PULSE(0 1.8 20m 0.1p 0.1p 20m 40m 200)
V12 d2 0 PULSE(0 1.8 40m 0.1p 0.1p 40m 80m 180)
V13 d3 0 PULSE(0 1.8 80m 0.1p 0.1p 80m 160m 150)
V14 d4 0 PULSE(0 1.8 160m 0.1p 0.1p 160m 320m 160)
V15 d5 0 PULSE(0 1.8 320m 0.1p 0.1p 320m 640m 80)

* block symbol definitions
.subckt 10bit d0 d1 d2 d3 d4 d5 d6 d7 d8 d9 10VrefIn Vo 10VrefOut
XX1 d0 d1 d2 d3 d4 d5 d6 d7 d8 10VrefIn N001 N002 9bit
XX2 d0 d1 d2 d3 d4 d5 d6 d7 d8 N002 N003 10VrefOut 9bit
XX3 d9 N001 N003 Vo switchbasic
.ends 10bit

.subckt 9bit d0 d1 d2 d3 d4 d5 d6 d7 d8 9VrefIn Vo 9VrefOut
XX1 d0 d1 d2 d3 d4 d5 d6 d7 9VrefIn N001 N002 8bit
XX2 d0 d1 d2 d3 d4 d5 d6 d7 N002 N003 9VrefOut 8bit
XX3 d8 N001 N003 Vo switchbasic
.ends 9bit

.subckt switchbasic d in_1 in_2 Vout
V1 N001 0 3.3
M5 Vout d_inv in_2 0 NMOS l=180n w=1.8u
M1 in_1 N002 Vout 0 NMOS l=180n w=1.8u
M2 d_inv d 0 0 NMOS l=180n w=1.8u
M3 Vout N002 in_2 Vout PMOS l=180n w=4u
M6 d_inv d N001 N001 PMOS l=180n w=4u
M7 Vout d_inv in_1 in_1 PMOS l=180n w=4u
M4 N002 d_inv 0 0 NMOS l=180n w=1.8u
M8 N002 d_inv N001 N001 PMOS l=180n w=1.8u
C1 Vout 0 1n
.ends switchbasic

.subckt 8bit d0 d1 d2 d3 d4 d5 d6 d7 8VrefIn Vo 8VrefOut
XX1 d0 d1 d2 d3 d4 d5 d6 8VrefIn N001 N003 7bit
XX2 d0 d1 d2 d3 d4 d5 d6 N003 N002 8VrefOut 7bit
XX3 d7 N001 N002 Vo switchbasic
.ends 8bit

.subckt 7bit d0 d1 d2 d3 d4 d5 d6 7VrefIn Vo 7VrefOut
XX1 d0 d1 d2 d3 d4 d5 7VrefIn N003 N001 6bit
XX2 d0 d1 d2 d3 d4 d5 N003 7VrefOut N002 6bit
XX3 d6 N001 N002 Vo switchbasic
.ends 7bit

.subckt 6bit d0 d1 d2 d3 d4 d5 6VrefIn 6VrefOut Vo
XX1 d0 d1 d2 d3 d4 6VrefIn N001 N002 5bit
XX2 d0 d1 d2 d3 d4 N002 N003 6VrefOut 5bit
XX3 d5 N001 N003 Vo switchbasic
.ends 6bit

.subckt 5bit d0 d1 d2 d3 d4 5VrefIn Vo 5VrefOut
XX1 d0 d1 d2 d3 5VrefIn N001 N002 4bit
XX2 d0 d1 d2 d3 N002 N003 5VrefOut 4bit
XX3 d4 N001 N003 Vo switchbasic
.ends 5bit

.subckt 4bit d0 d1 d2 d3 4VrefIn Vo 4VrefOut
XX1 d0 d1 d2 4VrefIn N001 N002 3bit
XX2 d0 d1 d2 N002 N003 4VrefOut 3bit
XX3 d3 N001 N003 Vo switchbasic
.ends 4bit

.subckt 3bit d0 d1 d2 3VrefIn Vo 3VrefOut
XX1 d0 d1 3VrefIn N002 N001 2bit
XX2 d0 d1 N002 3VrefOut N003 2bit
XX3 d2 N001 N003 Vo switchbasic
.ends 3bit

.subckt 2bit d0 d1 2VrefIn 2VrefOut Vo
XX1 d0 N001 N003 N002 switchbasic
R2 2VrefIn N001 100
R3 N001 N003 100
R4 N003 N005 100
XX2 d0 N005 2VrefOut N004 switchbasic
XX3 d1 N002 N004 Vo switchbasic
R1 N005 2VrefOut 100
.ends 2bit

.model NMOS NMOS (LEVEL=8 VERSION=3.2 TNOM=27 TOX=4.1E-9 XJ=1E-7 NCH=2.3549E17 VTH0=0.3823463 K1=0.5810697 
+            K2=4.774618E-3 K3=0.0431669 K3B=1.1498346 W0=1E-7 NLX=1.910552E-7 DVT0W=0 DVT1W=0 DVT2W=0 
+            DVT0=1.2894824 DVT1=0.3622063 DVT2=0.0713729 U0=280.633249 UA=-1.208537E-9 UB=2.158625E-18
+            UC=5.342807E-11 VSAT=9.366802E4 A0=1.7593146 AGS=0.3939741 B0=-6.413949E-9 B1=-1E-7 KETA=-5.180424E-4
+            A1=0 A2=1 RDSW=105.5517558 PRWG=0.5 PRWB=-0.1998871 WR=1 WINT=7.904732E-10 LINT=1.571424E-8 XL=0
+            XW=-1E-8 DWG=1.297221E-9 DWB=1.479041E-9 VOFF=-0.0955434 NFACTOR=2.4358891 CIT=0 CDSC=2.4E-4 CDSCD=0
+            CDSCB=0 ETA0=3.104851E-3 ETAB=-2.512384E-5 DSUB=0.0167075 PCLM=0.8073191 PDIBLC1=0.1666161 PDIBLC2=3.112892E-3    
+            PDIBLCB=-0.1 DROUT=0.7875618 PSCBE1=8E10 PSCBE2=9.213635E-10 PVAG=3.85243E-3 DELTA=0.01 RSH=6.7 MOBMOD=1
+            PRT=0 UTE=-1.5 KT1=-0.11 KT1L=0 KT2=0.022 UA1=4.31E-9 UB1=-7.61E-18 UC1=-5.6E-11 AT=3.3E4 WL=0 WLN=1
+            WW=0 WWN=1 WWL=0 LL=0 LLN=1 LW=0 LWN=1 LWL=0 CAPMOD=2 XPART=0.5 CGDO=7.08E-10 CGSO=7.08E-10 CGBO=1E-12
+            CJ=9.68858E-4 PB=0.8 MJ=0.3864502 CJSW=2.512138E-10 PBSW=0.809286 MJSW=0.1060414 CJSWG=3.3E-10 PBSWG=0.809286 
+            MJSWG=0.1060414 CF=0 PVTH0=-1.192722E-3 PRDSW=-5 PK2=6.450505E-5 WKETA=-4.27294E-4 LKETA=-0.0104078 
+            PU0=6.3268729 PUA=2.226552E-11 PUB=0 PVSAT=969.1480157 PETA0=1E-4 PKETA=-1.049509E-3)

.model PMOS PMOS (LEVEL=8 VERSION=3.2 TNOM=27 TOX=4.1E-9 XJ=1E-7 NCH=4.1589E17 VTH0=-0.3938813 K1=0.5479015
+            K2=0.0360586 K3=0.0993095 K3B=5.7086622 W0=1E-6 NLX=1.313191E-7 DVT0W=0 DVT1W=0 DVT2W=0 DVT0=0.4911363
+            DVT1=0.2227356 DVT2=0.1 U0=115.6852975 UA=1.505832E-9 UB=1E-21 UC=-1E-10 VSAT=1.329694E5 A0=1.7590478
+            AGS=0.3641621 B0=3.427126E-7 B1=1.062928E-6 KETA=0.0134667 A1=0.6859506 A2=0.3506788 RDSW=168.5705677
+            PRWG=0.5 PRWB=-0.4987371 WR=1 WINT=0 LINT=3.028832E-8 XL=0 XW=-1E-8 DWG=-2.349633E-8 DWB=-7.152486E-9 
+            VOFF=-0.0994037 NFACTOR=1.9424315 CIT=0 CDSC=2.4E-4 CDSCD=0 CDSCB=0 ETA0=0.0608072 ETAB=-0.0426148
+            DSUB=0.7343015 PCLM=3.2579974 PDIBLC1=7.229527E-6 PDIBLC2=0.025389 PDIBLCB=-1E-3 DROUT=0 PSCBE1=1.454878E10
+            PSCBE2=4.202027E-9 PVAG=15 DELTA=0.01 RSH=7.8 MOBMOD=1 PRT=0 UTE=-1.5 KT1=-0.11 KT1L=0 KT2=0.022 UA1=4.31E-9
+            UB1=-7.61E-18 UC1=-5.6E-11 AT=3.3E4 WL=0 WLN=1 WW=0 WWN=1 WWL=0 LL=0 LLN=1 LW=0 LWN=1 LWL=0 CAPMOD=2 XPART=0.5
+            CGDO=6.32E-10 CGSO=6.32E-10 CGBO=1E-12 CJ=1.172138E-3 PB=0.8421173 MJ=0.4109788 CJSW=2.242609E-10 PBSW=0.8            
+            MJSW=0.3752089 CJSWG=4.22E-10 PBSWG=0.8 MJSWG=0.3752089 CF=0 PVTH0=1.888482E-3 PRDSW=11.5315407 PK2=1.559399E-3    
+            WKETA=0.0319301 LKETA=2.955547E-3 PU0=-1.1105313 PUA=-4.62102E-11 PUB=1E-21 PVSAT=50 PETA0=1E-4 PKETA=-4.346368E-3)

.tran 10ms 10s
.control
run
plot v(out)
.endc
.end
